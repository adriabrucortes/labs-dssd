`include "../misc/timescale.v"

module tb_top_meteo_de0cv();

  TO BE COMPLETED BY THE STUDENT

endmodule
